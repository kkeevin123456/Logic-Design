module MO(clk, reset, in_data, i, j, opcode, out_data, fin);
input clk, reset;
input [9:0] in_data;
output fin;
output [2:0] opcode;
output [9:0] i, j;
output [19:0] out_data;

//(your code)...

endmodule